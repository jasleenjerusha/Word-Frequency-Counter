
module counter ( clk, reset, enable, dat_out );
  output [15:0] dat_out;
  input clk, reset, enable;
  wire   N69, N70, N71, N72, N73, N74, N75, N76, N77, N78, N79, N80, N81, N82,
         N83, N84, N86, N88, N90, N92, N94, N96, n42, n43, n44, n45, n46, n47,
         n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61,
         n62, n63, n64, n65, n66, n67;

endmodule

///////////////

module submod (in1, in2, out1);
 output out1;
 input in1, in2;

wire N01;

endmodule

//////////////

module submod1 (in1, in2, out1);
 output out1;
 input in1, in2;

wire N01;

endmodule

